library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package dtype_memc_ord_pkg is
    type t_cmp_ord is record
{pkg_signals}
    end record t_cmp_ord;
end package;